// Code your design here
`include "struct_diag.sv"
`include "alarm.sv"
`include "ct_mod_N.sv"
`include "lcd_int3.sv"